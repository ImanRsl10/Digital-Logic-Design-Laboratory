library verilog;
use verilog.vl_types.all;
entity Wrapper_TB is
end Wrapper_TB;
