library verilog;
use verilog.vl_types.all;
entity Wrapper_PostSynthesis_TB is
end Wrapper_PostSynthesis_TB;
